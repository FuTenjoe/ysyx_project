`include "../vsrc/rvseed_defines.v"

module clint  (
/*    input clk,
    input rst_n*/
);
    




endmodule
`include "../vsrc/rvseed_defines.v"

module cache_axi_judge (
    input mem_req,
    input mem_valid
);


endmodule
`include "../vsrc/rvseed_defines.v"

module cache_axi_judge (
    input if_valid,
    input waxi_valid,
    input w_done,
    input dd_r_done2,
    output cpu_req
);


endmodule